
module and_gate (
  input a,  
  input b,
  output q
);

assign q = a && b;

endmodule
